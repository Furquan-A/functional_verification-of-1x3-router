class wr_agt_config extends uvm_object;
`uvm_object_utils(wr_agt_config)

bit has_monitor = 1;
bit 