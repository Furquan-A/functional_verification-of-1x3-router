class wr_driver extends uvm_driver;
`uvm_component_utils(wr_driver)

wr_agt_config m_cfg;